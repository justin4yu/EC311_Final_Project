module bcd_converter(

);

endmodule;